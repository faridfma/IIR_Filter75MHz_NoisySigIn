library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


-- this codde use DSS to test Butterworth IIR fillter
--Fs = 1.55MHz; Fpass=37.5Khz, Fstop = 200KHz; Astop = 40dB; Apass = 1dB

entity IIR_Filter_Pipelined_ChbyChevII_Fc37K5_Fp100K_Astop60Test is
    Port (
        clk                  : in  std_logic := '0';           -- Clock signal
        ce                   : in  std_logic := '0'; 
        reset                : in  std_logic := '0';           -- Reset signal
      --  x_in                 : in  std_logic_vector(15 downto 0):= (others=>'0');  -- Input signal x[n] (Q0.16 format) 
        x_in                 : in  signed (15 downto 0):= (others=>'0');  -- Input signal x[n] (Q0.16 format)
        --x_in_out             : Out std_logic_vector(15 downto 0):= (others=>'0');   
        iir_out              : out std_logic_vector(15 downto 0):= (others=>'0');  -- Filtered output
        sample_valid_in      : out std_logic := '0';      -- Sample valid input signal
        sample_valid_out     : out std_logic := '0';     -- Sample valid output signal
        busy                 : out std_logic := '0'      -- Busy signal
    );
end IIR_Filter_Pipelined_ChbyChevII_Fc37K5_Fp100K_Astop60Test;

architecture Behavioral of IIR_Filter_Pipelined_ChbyChevII_Fc37K5_Fp100K_Astop60Test is


    signal x_in_Sig : signed (15 downto 0):= (others=>'0');  -- Input signal x[n] (Q0.16 format)
 
    -- Register declarations for input (x) and output (y) values
    type x_regArray is array(0 to 6) of signed(31 downto 0);  -- Input registers (x); add 8 bits for scaling
    signal x_reg : x_regArray; 
    type y_regArray is array(0 to 6) of signed(31 downto 0);  -- Input registers (y)
    signal y_reg : y_regArray; 

    -- Multiplication signals
   type mul_xArray  is array(0 to 6) of signed(63 downto 0); --16 bits times 8 bits ==>24 bits
   signal mul_x : mul_xArray; 
   type mul_yArray is array(1 to 6) of signed(63 downto 0);  --16 bits times 8 bits ==>24 bits
   signal mul_y : mul_yArray; 
   
   -- Sum signals
   type Sum_xArray is array(0 to 6) of signed(63 downto 0);  -- need 27 bits
   signal Sum_x : Sum_xArray;  
   type Sum_yArray  is array(0 to 6) of signed(63 downto 0);  --need 26 bits
   signal Sum_y : Sum_yArray; 
    
   -- Coefficients (b and a arrays)
   type b_Coefficients is array(0 to 6) of signed(31 downto 0);
   type a_Coefficients is array(0 to 6) of signed(31 downto 0);
    
   constant b : b_Coefficients := (
--        to_signed(15, 32),
--        to_signed(61, 32),
--        to_signed(91, 32),
--        to_signed(61, 32),
--        to_signed(15, 32)
        
        to_signed(20004, 32),
        to_signed(-79756, 32),
        to_signed(154737, 32),
        to_signed(-188354, 32),
        to_signed(154737, 32),
        to_signed(-79756, 32),
        to_signed(20004, 32)       
    );

    constant a : a_Coefficients := (
--        to_signed(65536, 32),
--        to_signed(-216338, 32),
--        to_signed(271135, 32),
--        to_signed(-152556, 32),
--        to_signed(32466, 32)
        
        to_signed(16777216, 32),
        to_signed(-86221058, 32),
        to_signed(185542407, 32),
        to_signed(-213901648, 32),
        to_signed(139278978, 32),
        to_signed(-48550822, 32),
        to_signed(7076543, 32)

    );
    

    -- Final output signal
    signal Output : signed(31 downto 0):= (others=>'0');  
    
    signal OutputX : signed(63 downto 0):= (others=>'0'); 
    signal OutputY : signed(63 downto 0):= (others=>'0'); 

    -- State machine state
    signal state : integer := 0;


    signal sample_validin_Sig: std_logic := '0'; 
    signal clockcounter : integer range 0 to 64;  

    signal Flag: std_logic := '0'; 

    type InputData_Array is array(0 to 1559) of signed(15 downto 0);  -- need 27 bits
    signal InputData : InputData_Array := (  
    
    to_signed(0,16),
    to_signed(8160,16),
    to_signed(-9127,16),
    to_signed(11676,16),
    to_signed(894,16),
    to_signed(-710,16),
    to_signed(15512,16),
    to_signed(-4154,16),
    to_signed(12049,16),
    to_signed(10408,16),
    to_signed(-428,16),
    to_signed(20301,16),
    to_signed(2922,16),
    to_signed(10973,16),
    to_signed(19005,16),
    to_signed(1574,16),
    to_signed(22214,16),
    to_signed(11253,16),
    to_signed(9453,16),
    to_signed(25462,16),
    to_signed(5567,16),
    to_signed(21526,16),
    to_signed(19625,16),
    to_signed(8514,16),
    to_signed(28953,16),
    to_signed(11272,16),
    to_signed(19005,16),
    to_signed(26708,16),
    to_signed(8934,16),
    to_signed(29220,16),
    to_signed(17893,16),
    to_signed(15717,16),
    to_signed(31339,16),
    to_signed(11048,16),
    to_signed(26601,16),
    to_signed(24287,16),
    to_signed(12755,16),
    to_signed(32767,16),
    to_signed(14651,16),
    to_signed(21945,16),
    to_signed(29204,16),
    to_signed(10982,16),
    to_signed(30816,16),
    to_signed(19035,16),
    to_signed(16403,16),
    to_signed(31567,16),
    to_signed(10819,16),
    to_signed(25915,16),
    to_signed(23145,16),
    to_signed(11159,16),
    to_signed(30719,16),
    to_signed(12155,16),
    to_signed(19005,16),
    to_signed(25824,16),
    to_signed(7168,16),
    to_signed(26574,16),
    to_signed(14373,16),
    to_signed(11327,16),
    to_signed(26087,16),
    to_signed(4942,16),
    to_signed(19652,16),
    to_signed(16505,16),
    to_signed(4153,16),
    to_signed(23359,16),
    to_signed(4453,16),
    to_signed(10973,16),
    to_signed(17475,16),
    to_signed(-1485,16),
    to_signed(17632,16),
    to_signed(5156,16),
    to_signed(1850,16),
    to_signed(16365,16),
    to_signed(-5008,16),
    to_signed(9489,16),
    to_signed(6146,16),
    to_signed(-6385,16),
    to_signed(12659,16),
    to_signed(-6393,16),
    to_signed(0,16),
    to_signed(6393,16),
    to_signed(-12659,16),
    to_signed(6385,16),
    to_signed(-6146,16),
    to_signed(-9489,16),
    to_signed(5008,16),
    to_signed(-16365,16),
    to_signed(-1850,16),
    to_signed(-5156,16),
    to_signed(-17632,16),
    to_signed(1485,16),
    to_signed(-17475,16),
    to_signed(-10973,16),
    to_signed(-4453,16),
    to_signed(-23359,16),
    to_signed(-4153,16),
    to_signed(-16505,16),
    to_signed(-19652,16),
    to_signed(-4942,16),
    to_signed(-26087,16),
    to_signed(-11327,16),
    to_signed(-14373,16),
    to_signed(-26574,16),
    to_signed(-7168,16),
    to_signed(-25824,16),
    to_signed(-19005,16),
    to_signed(-12155,16),
    to_signed(-30719,16),
    to_signed(-11159,16),
    to_signed(-23145,16),
    to_signed(-25915,16),
    to_signed(-10819,16),
    to_signed(-31567,16),
    to_signed(-16403,16),
    to_signed(-19035,16),
    to_signed(-30816,16),
    to_signed(-10982,16),
    to_signed(-29204,16),
    to_signed(-21945,16),
    to_signed(-14651,16),
    to_signed(-32767,16),
    to_signed(-12755,16),
    to_signed(-24287,16),
    to_signed(-26601,16),
    to_signed(-11048,16),
    to_signed(-31339,16),
    to_signed(-15717,16),
    to_signed(-17893,16),
    to_signed(-29220,16),
    to_signed(-8934,16),
    to_signed(-26708,16),
    to_signed(-19005,16),
    to_signed(-11272,16),
    to_signed(-28953,16),
    to_signed(-8514,16),
    to_signed(-19625,16),
    to_signed(-21526,16),
    to_signed(-5567,16),
    to_signed(-25462,16),
    to_signed(-9453,16),
    to_signed(-11253,16),
    to_signed(-22214,16),
    to_signed(-1574,16),
    to_signed(-19005,16),
    to_signed(-10973,16),
    to_signed(-2922,16),
    to_signed(-20301,16),
    to_signed(428,16),
    to_signed(-10408,16),
    to_signed(-12049,16),
    to_signed(4154,16),
    to_signed(-15512,16),
    to_signed(710,16),
    to_signed(-894,16),
    to_signed(-11676,16),
    to_signed(9127,16),
    to_signed(-8160,16),
    to_signed(0,16),
    to_signed(8160,16),
    to_signed(-9127,16),
    to_signed(11676,16),
    to_signed(894,16),
    to_signed(-710,16),
    to_signed(15512,16),
    to_signed(-4154,16),
    to_signed(12049,16),
    to_signed(10408,16),
    to_signed(-428,16),
    to_signed(20301,16),
    to_signed(2922,16),
    to_signed(10973,16),
    to_signed(19005,16),
    to_signed(1574,16),
    to_signed(22214,16),
    to_signed(11253,16),
    to_signed(9453,16),
    to_signed(25462,16),
    to_signed(5567,16),
    to_signed(21526,16),
    to_signed(19625,16),
    to_signed(8514,16),
    to_signed(28953,16),
    to_signed(11272,16),
    to_signed(19005,16),
    to_signed(26708,16),
    to_signed(8934,16),
    to_signed(29220,16),
    to_signed(17893,16),
    to_signed(15717,16),
    to_signed(31339,16),
    to_signed(11048,16),
    to_signed(26601,16),
    to_signed(24287,16),
    to_signed(12755,16),
    to_signed(32767,16),
    to_signed(14651,16),
    to_signed(21945,16),
    to_signed(29204,16),
    to_signed(10982,16),
    to_signed(30816,16),
    to_signed(19035,16),
    to_signed(16403,16),
    to_signed(31567,16),
    to_signed(10819,16),
    to_signed(25915,16),
    to_signed(23145,16),
    to_signed(11159,16),
    to_signed(30719,16),
    to_signed(12155,16),
    to_signed(19005,16),
    to_signed(25824,16),
    to_signed(7168,16),
    to_signed(26574,16),
    to_signed(14373,16),
    to_signed(11327,16),
    to_signed(26087,16),
    to_signed(4942,16),
    to_signed(19652,16),
    to_signed(16505,16),
    to_signed(4153,16),
    to_signed(23359,16),
    to_signed(4453,16),
    to_signed(10973,16),
    to_signed(17475,16),
    to_signed(-1485,16),
    to_signed(17632,16),
    to_signed(5156,16),
    to_signed(1850,16),
    to_signed(16365,16),
    to_signed(-5008,16),
    to_signed(9489,16),
    to_signed(6146,16),
    to_signed(-6385,16),
    to_signed(12659,16),
    to_signed(-6393,16),
    to_signed(0,16),
    to_signed(6393,16),
    to_signed(-12659,16),
    to_signed(6385,16),
    to_signed(-6146,16),
    to_signed(-9489,16),
    to_signed(5008,16),
    to_signed(-16365,16),
    to_signed(-1850,16),
    to_signed(-5156,16),
    to_signed(-17632,16),
    to_signed(1485,16),
    to_signed(-17475,16),
    to_signed(-10973,16),
    to_signed(-4453,16),
    to_signed(-23359,16),
    to_signed(-4153,16),
    to_signed(-16505,16),
    to_signed(-19652,16),
    to_signed(-4942,16),
    to_signed(-26087,16),
    to_signed(-11327,16),
    to_signed(-14373,16),
    to_signed(-26574,16),
    to_signed(-7168,16),
    to_signed(-25824,16),
    to_signed(-19005,16),
    to_signed(-12155,16),
    to_signed(-30719,16),
    to_signed(-11159,16),
    to_signed(-23145,16),
    to_signed(-25915,16),
    to_signed(-10819,16),
    to_signed(-31567,16),
    to_signed(-16403,16),
    to_signed(-19035,16),
    to_signed(-30816,16),
    to_signed(-10982,16),
    to_signed(-29204,16),
    to_signed(-21945,16),
    to_signed(-14651,16),
    to_signed(-32767,16),
    to_signed(-12755,16),
    to_signed(-24287,16),
    to_signed(-26601,16),
    to_signed(-11048,16),
    to_signed(-31339,16),
    to_signed(-15717,16),
    to_signed(-17893,16),
    to_signed(-29220,16),
    to_signed(-8934,16),
    to_signed(-26708,16),
    to_signed(-19005,16),
    to_signed(-11272,16),
    to_signed(-28953,16),
    to_signed(-8514,16),
    to_signed(-19625,16),
    to_signed(-21526,16),
    to_signed(-5567,16),
    to_signed(-25462,16),
    to_signed(-9453,16),
    to_signed(-11253,16),
    to_signed(-22214,16),
    to_signed(-1574,16),
    to_signed(-19005,16),
    to_signed(-10973,16),
    to_signed(-2922,16),
    to_signed(-20301,16),
    to_signed(428,16),
    to_signed(-10408,16),
    to_signed(-12049,16),
    to_signed(4154,16),
    to_signed(-15512,16),
    to_signed(710,16),
    to_signed(-894,16),
    to_signed(-11676,16),
    to_signed(9127,16),
    to_signed(-8160,16),
    to_signed(0,16),
    to_signed(8160,16),
    to_signed(-9127,16),
    to_signed(11676,16),
    to_signed(894,16),
    to_signed(-710,16),
    to_signed(15512,16),
    to_signed(-4154,16),
    to_signed(12049,16),
    to_signed(10408,16),
    to_signed(-428,16),
    to_signed(20301,16),
    to_signed(2922,16),
    to_signed(10973,16),
    to_signed(19005,16),
    to_signed(1574,16),
    to_signed(22214,16),
    to_signed(11253,16),
    to_signed(9453,16),
    to_signed(25462,16),
    to_signed(5567,16),
    to_signed(21526,16),
    to_signed(19625,16),
    to_signed(8514,16),
    to_signed(28953,16),
    to_signed(11272,16),
    to_signed(19005,16),
    to_signed(26708,16),
    to_signed(8934,16),
    to_signed(29220,16),
    to_signed(17893,16),
    to_signed(15717,16),
    to_signed(31339,16),
    to_signed(11048,16),
    to_signed(26601,16),
    to_signed(24287,16),
    to_signed(12755,16),
    to_signed(32767,16),
    to_signed(14651,16),
    to_signed(21945,16),
    to_signed(29204,16),
    to_signed(10982,16),
    to_signed(30816,16),
    to_signed(19035,16),
    to_signed(16403,16),
    to_signed(31567,16),
    to_signed(10819,16),
    to_signed(25915,16),
    to_signed(23145,16),
    to_signed(11159,16),
    to_signed(30719,16),
    to_signed(12155,16),
    to_signed(19005,16),
    to_signed(25824,16),
    to_signed(7168,16),
    to_signed(26574,16),
    to_signed(14373,16),
    to_signed(11327,16),
    to_signed(26087,16),
    to_signed(4942,16),
    to_signed(19652,16),
    to_signed(16505,16),
    to_signed(4153,16),
    to_signed(23359,16),
    to_signed(4453,16),
    to_signed(10973,16),
    to_signed(17475,16),
    to_signed(-1485,16),
    to_signed(17632,16),
    to_signed(5156,16),
    to_signed(1850,16),
    to_signed(16365,16),
    to_signed(-5008,16),
    to_signed(9489,16),
    to_signed(6146,16),
    to_signed(-6385,16),
    to_signed(12659,16),
    to_signed(-6393,16),
    to_signed(0,16),
    to_signed(6393,16),
    to_signed(-12659,16),
    to_signed(6385,16),
    to_signed(-6146,16),
    to_signed(-9489,16),
    to_signed(5008,16),
    to_signed(-16365,16),
    to_signed(-1850,16),
    to_signed(-5156,16),
    to_signed(-17632,16),
    to_signed(1485,16),
    to_signed(-17475,16),
    to_signed(-10973,16),
    to_signed(-4453,16),
    to_signed(-23359,16),
    to_signed(-4153,16),
    to_signed(-16505,16),
    to_signed(-19652,16),
    to_signed(-4942,16),
    to_signed(-26087,16),
    to_signed(-11327,16),
    to_signed(-14373,16),
    to_signed(-26574,16),
    to_signed(-7168,16),
    to_signed(-25824,16),
    to_signed(-19005,16),
    to_signed(-12155,16),
    to_signed(-30719,16),
    to_signed(-11159,16),
    to_signed(-23145,16),
    to_signed(-25915,16),
    to_signed(-10819,16),
    to_signed(-31567,16),
    to_signed(-16403,16),
    to_signed(-19035,16),
    to_signed(-30816,16),
    to_signed(-10982,16),
    to_signed(-29204,16),
    to_signed(-21945,16),
    to_signed(-14651,16),
    to_signed(-32767,16),
    to_signed(-12755,16),
    to_signed(-24287,16),
    to_signed(-26601,16),
    to_signed(-11048,16),
    to_signed(-31339,16),
    to_signed(-15717,16),
    to_signed(-17893,16),
    to_signed(-29220,16),
    to_signed(-8934,16),
    to_signed(-26708,16),
    to_signed(-19005,16),
    to_signed(-11272,16),
    to_signed(-28953,16),
    to_signed(-8514,16),
    to_signed(-19625,16),
    to_signed(-21526,16),
    to_signed(-5567,16),
    to_signed(-25462,16),
    to_signed(-9453,16),
    to_signed(-11253,16),
    to_signed(-22214,16),
    to_signed(-1574,16),
    to_signed(-19005,16),
    to_signed(-10973,16),
    to_signed(-2922,16),
    to_signed(-20301,16),
    to_signed(428,16),
    to_signed(-10408,16),
    to_signed(-12049,16),
    to_signed(4154,16),
    to_signed(-15512,16),
    to_signed(710,16),
    to_signed(-894,16),
    to_signed(-11676,16),
    to_signed(9127,16),
    to_signed(-8160,16),
    to_signed(0,16),
    to_signed(8160,16),
    to_signed(-9127,16),
    to_signed(11676,16),
    to_signed(894,16),
    to_signed(-710,16),
    to_signed(15512,16),
    to_signed(-4154,16),
    to_signed(12049,16),
    to_signed(10408,16),
    to_signed(-428,16),
    to_signed(20301,16),
    to_signed(2922,16),
    to_signed(10973,16),
    to_signed(19005,16),
    to_signed(1574,16),
    to_signed(22214,16),
    to_signed(11253,16),
    to_signed(9453,16),
    to_signed(25462,16),
    to_signed(5567,16),
    to_signed(21526,16),
    to_signed(19625,16),
    to_signed(8514,16),
    to_signed(28953,16),
    to_signed(11272,16),
    to_signed(19005,16),
    to_signed(26708,16),
    to_signed(8934,16),
    to_signed(29220,16),
    to_signed(17893,16),
    to_signed(15717,16),
    to_signed(31339,16),
    to_signed(11048,16),
    to_signed(26601,16),
    to_signed(24287,16),
    to_signed(12755,16),
    to_signed(32767,16),
    to_signed(14651,16),
    to_signed(21945,16),
    to_signed(29204,16),
    to_signed(10982,16),
    to_signed(30816,16),
    to_signed(19035,16),
    to_signed(16403,16),
    to_signed(31567,16),
    to_signed(10819,16),
    to_signed(25915,16),
    to_signed(23145,16),
    to_signed(11159,16),
    to_signed(30719,16),
    to_signed(12155,16),
    to_signed(19005,16),
    to_signed(25824,16),
    to_signed(7168,16),
    to_signed(26574,16),
    to_signed(14373,16),
    to_signed(11327,16),
    to_signed(26087,16),
    to_signed(4942,16),
    to_signed(19652,16),
    to_signed(16505,16),
    to_signed(4153,16),
    to_signed(23359,16),
    to_signed(4453,16),
    to_signed(10973,16),
    to_signed(17475,16),
    to_signed(-1485,16),
    to_signed(17632,16),
    to_signed(5156,16),
    to_signed(1850,16),
    to_signed(16365,16),
    to_signed(-5008,16),
    to_signed(9489,16),
    to_signed(6146,16),
    to_signed(-6385,16),
    to_signed(12659,16),
    to_signed(-6393,16),
    to_signed(0,16),
    to_signed(6393,16),
    to_signed(-12659,16),
    to_signed(6385,16),
    to_signed(-6146,16),
    to_signed(-9489,16),
    to_signed(5008,16),
    to_signed(-16365,16),
    to_signed(-1850,16),
    to_signed(-5156,16),
    to_signed(-17632,16),
    to_signed(1485,16),
    to_signed(-17475,16),
    to_signed(-10973,16),
    to_signed(-4453,16),
    to_signed(-23359,16),
    to_signed(-4153,16),
    to_signed(-16505,16),
    to_signed(-19652,16),
    to_signed(-4942,16),
    to_signed(-26087,16),
    to_signed(-11327,16),
    to_signed(-14373,16),
    to_signed(-26574,16),
    to_signed(-7168,16),
    to_signed(-25824,16),
    to_signed(-19005,16),
    to_signed(-12155,16),
    to_signed(-30719,16),
    to_signed(-11159,16),
    to_signed(-23145,16),
    to_signed(-25915,16),
    to_signed(-10819,16),
    to_signed(-31567,16),
    to_signed(-16403,16),
    to_signed(-19035,16),
    to_signed(-30816,16),
    to_signed(-10982,16),
    to_signed(-29204,16),
    to_signed(-21945,16),
    to_signed(-14651,16),
    to_signed(-32767,16),
    to_signed(-12755,16),
    to_signed(-24287,16),
    to_signed(-26601,16),
    to_signed(-11048,16),
    to_signed(-31339,16),
    to_signed(-15717,16),
    to_signed(-17893,16),
    to_signed(-29220,16),
    to_signed(-8934,16),
    to_signed(-26708,16),
    to_signed(-19005,16),
    to_signed(-11272,16),
    to_signed(-28953,16),
    to_signed(-8514,16),
    to_signed(-19625,16),
    to_signed(-21526,16),
    to_signed(-5567,16),
    to_signed(-25462,16),
    to_signed(-9453,16),
    to_signed(-11253,16),
    to_signed(-22214,16),
    to_signed(-1574,16),
    to_signed(-19005,16),
    to_signed(-10973,16),
    to_signed(-2922,16),
    to_signed(-20301,16),
    to_signed(428,16),
    to_signed(-10408,16),
    to_signed(-12049,16),
    to_signed(4154,16),
    to_signed(-15512,16),
    to_signed(710,16),
    to_signed(-894,16),
    to_signed(-11676,16),
    to_signed(9127,16),
    to_signed(-8160,16),
    to_signed(0,16),
    to_signed(8160,16),
    to_signed(-9127,16),
    to_signed(11676,16),
    to_signed(894,16),
    to_signed(-710,16),
    to_signed(15512,16),
    to_signed(-4154,16),
    to_signed(12049,16),
    to_signed(10408,16),
    to_signed(-428,16),
    to_signed(20301,16),
    to_signed(2922,16),
    to_signed(10973,16),
    to_signed(19005,16),
    to_signed(1574,16),
    to_signed(22214,16),
    to_signed(11253,16),
    to_signed(9453,16),
    to_signed(25462,16),
    to_signed(5567,16),
    to_signed(21526,16),
    to_signed(19625,16),
    to_signed(8514,16),
    to_signed(28953,16),
    to_signed(11272,16),
    to_signed(19005,16),
    to_signed(26708,16),
    to_signed(8934,16),
    to_signed(29220,16),
    to_signed(17893,16),
    to_signed(15717,16),
    to_signed(31339,16),
    to_signed(11048,16),
    to_signed(26601,16),
    to_signed(24287,16),
    to_signed(12755,16),
    to_signed(32767,16),
    to_signed(14651,16),
    to_signed(21945,16),
    to_signed(29204,16),
    to_signed(10982,16),
    to_signed(30816,16),
    to_signed(19035,16),
    to_signed(16403,16),
    to_signed(31567,16),
    to_signed(10819,16),
    to_signed(25915,16),
    to_signed(23145,16),
    to_signed(11159,16),
    to_signed(30719,16),
    to_signed(12155,16),
    to_signed(19005,16),
    to_signed(25824,16),
    to_signed(7168,16),
    to_signed(26574,16),
    to_signed(14373,16),
    to_signed(11327,16),
    to_signed(26087,16),
    to_signed(4942,16),
    to_signed(19652,16),
    to_signed(16505,16),
    to_signed(4153,16),
    to_signed(23359,16),
    to_signed(4453,16),
    to_signed(10973,16),
    to_signed(17475,16),
    to_signed(-1485,16),
    to_signed(17632,16),
    to_signed(5156,16),
    to_signed(1850,16),
    to_signed(16365,16),
    to_signed(-5008,16),
    to_signed(9489,16),
    to_signed(6146,16),
    to_signed(-6385,16),
    to_signed(12659,16),
    to_signed(-6393,16),
    to_signed(0,16),
    to_signed(6393,16),
    to_signed(-12659,16),
    to_signed(6385,16),
    to_signed(-6146,16),
    to_signed(-9489,16),
    to_signed(5008,16),
    to_signed(-16365,16),
    to_signed(-1850,16),
    to_signed(-5156,16),
    to_signed(-17632,16),
    to_signed(1485,16),
    to_signed(-17475,16),
    to_signed(-10973,16),
    to_signed(-4453,16),
    to_signed(-23359,16),
    to_signed(-4153,16),
    to_signed(-16505,16),
    to_signed(-19652,16),
    to_signed(-4942,16),
    to_signed(-26087,16),
    to_signed(-11327,16),
    to_signed(-14373,16),
    to_signed(-26574,16),
    to_signed(-7168,16),
    to_signed(-25824,16),
    to_signed(-19005,16),
    to_signed(-12155,16),
    to_signed(-30719,16),
    to_signed(-11159,16),
    to_signed(-23145,16),
    to_signed(-25915,16),
    to_signed(-10819,16),
    to_signed(-31567,16),
    to_signed(-16403,16),
    to_signed(-19035,16),
    to_signed(-30816,16),
    to_signed(-10982,16),
    to_signed(-29204,16),
    to_signed(-21945,16),
    to_signed(-14651,16),
    to_signed(-32767,16),
    to_signed(-12755,16),
    to_signed(-24287,16),
    to_signed(-26601,16),
    to_signed(-11048,16),
    to_signed(-31339,16),
    to_signed(-15717,16),
    to_signed(-17893,16),
    to_signed(-29220,16),
    to_signed(-8934,16),
    to_signed(-26708,16),
    to_signed(-19005,16),
    to_signed(-11272,16),
    to_signed(-28953,16),
    to_signed(-8514,16),
    to_signed(-19625,16),
    to_signed(-21526,16),
    to_signed(-5567,16),
    to_signed(-25462,16),
    to_signed(-9453,16),
    to_signed(-11253,16),
    to_signed(-22214,16),
    to_signed(-1574,16),
    to_signed(-19005,16),
    to_signed(-10973,16),
    to_signed(-2922,16),
    to_signed(-20301,16),
    to_signed(428,16),
    to_signed(-10408,16),
    to_signed(-12049,16),
    to_signed(4154,16),
    to_signed(-15512,16),
    to_signed(710,16),
    to_signed(-894,16),
    to_signed(-11676,16),
    to_signed(9127,16),
    to_signed(-8160,16),
    to_signed(0,16),
    to_signed(8160,16),
    to_signed(-9127,16),
    to_signed(11676,16),
    to_signed(894,16),
    to_signed(-710,16),
    to_signed(15512,16),
    to_signed(-4154,16),
    to_signed(12049,16),
    to_signed(10408,16),
    to_signed(-428,16),
    to_signed(20301,16),
    to_signed(2922,16),
    to_signed(10973,16),
    to_signed(19005,16),
    to_signed(1574,16),
    to_signed(22214,16),
    to_signed(11253,16),
    to_signed(9453,16),
    to_signed(25462,16),
    to_signed(5567,16),
    to_signed(21526,16),
    to_signed(19625,16),
    to_signed(8514,16),
    to_signed(28953,16),
    to_signed(11272,16),
    to_signed(19005,16),
    to_signed(26708,16),
    to_signed(8934,16),
    to_signed(29220,16),
    to_signed(17893,16),
    to_signed(15717,16),
    to_signed(31339,16),
    to_signed(11048,16),
    to_signed(26601,16),
    to_signed(24287,16),
    to_signed(12755,16),
    to_signed(32767,16),
    to_signed(14651,16),
    to_signed(21945,16),
    to_signed(29204,16),
    to_signed(10982,16),
    to_signed(30816,16),
    to_signed(19035,16),
    to_signed(16403,16),
    to_signed(31567,16),
    to_signed(10819,16),
    to_signed(25915,16),
    to_signed(23145,16),
    to_signed(11159,16),
    to_signed(30719,16),
    to_signed(12155,16),
    to_signed(19005,16),
    to_signed(25824,16),
    to_signed(7168,16),
    to_signed(26574,16),
    to_signed(14373,16),
    to_signed(11327,16),
    to_signed(26087,16),
    to_signed(4942,16),
    to_signed(19652,16),
    to_signed(16505,16),
    to_signed(4153,16),
    to_signed(23359,16),
    to_signed(4453,16),
    to_signed(10973,16),
    to_signed(17475,16),
    to_signed(-1485,16),
    to_signed(17632,16),
    to_signed(5156,16),
    to_signed(1850,16),
    to_signed(16365,16),
    to_signed(-5008,16),
    to_signed(9489,16),
    to_signed(6146,16),
    to_signed(-6385,16),
    to_signed(12659,16),
    to_signed(-6393,16),
    to_signed(0,16),
    to_signed(6393,16),
    to_signed(-12659,16),
    to_signed(6385,16),
    to_signed(-6146,16),
    to_signed(-9489,16),
    to_signed(5008,16),
    to_signed(-16365,16),
    to_signed(-1850,16),
    to_signed(-5156,16),
    to_signed(-17632,16),
    to_signed(1485,16),
    to_signed(-17475,16),
    to_signed(-10973,16),
    to_signed(-4453,16),
    to_signed(-23359,16),
    to_signed(-4153,16),
    to_signed(-16505,16),
    to_signed(-19652,16),
    to_signed(-4942,16),
    to_signed(-26087,16),
    to_signed(-11327,16),
    to_signed(-14373,16),
    to_signed(-26574,16),
    to_signed(-7168,16),
    to_signed(-25824,16),
    to_signed(-19005,16),
    to_signed(-12155,16),
    to_signed(-30719,16),
    to_signed(-11159,16),
    to_signed(-23145,16),
    to_signed(-25915,16),
    to_signed(-10819,16),
    to_signed(-31567,16),
    to_signed(-16403,16),
    to_signed(-19035,16),
    to_signed(-30816,16),
    to_signed(-10982,16),
    to_signed(-29204,16),
    to_signed(-21945,16),
    to_signed(-14651,16),
    to_signed(-32767,16),
    to_signed(-12755,16),
    to_signed(-24287,16),
    to_signed(-26601,16),
    to_signed(-11048,16),
    to_signed(-31339,16),
    to_signed(-15717,16),
    to_signed(-17893,16),
    to_signed(-29220,16),
    to_signed(-8934,16),
    to_signed(-26708,16),
    to_signed(-19005,16),
    to_signed(-11272,16),
    to_signed(-28953,16),
    to_signed(-8514,16),
    to_signed(-19625,16),
    to_signed(-21526,16),
    to_signed(-5567,16),
    to_signed(-25462,16),
    to_signed(-9453,16),
    to_signed(-11253,16),
    to_signed(-22214,16),
    to_signed(-1574,16),
    to_signed(-19005,16),
    to_signed(-10973,16),
    to_signed(-2922,16),
    to_signed(-20301,16),
    to_signed(428,16),
    to_signed(-10408,16),
    to_signed(-12049,16),
    to_signed(4154,16),
    to_signed(-15512,16),
    to_signed(710,16),
    to_signed(-894,16),
    to_signed(-11676,16),
    to_signed(9127,16),
    to_signed(-8160,16),
    to_signed(0,16),
    to_signed(8160,16),
    to_signed(-9127,16),
    to_signed(11676,16),
    to_signed(894,16),
    to_signed(-710,16),
    to_signed(15512,16),
    to_signed(-4154,16),
    to_signed(12049,16),
    to_signed(10408,16),
    to_signed(-428,16),
    to_signed(20301,16),
    to_signed(2922,16),
    to_signed(10973,16),
    to_signed(19005,16),
    to_signed(1574,16),
    to_signed(22214,16),
    to_signed(11253,16),
    to_signed(9453,16),
    to_signed(25462,16),
    to_signed(5567,16),
    to_signed(21526,16),
    to_signed(19625,16),
    to_signed(8514,16),
    to_signed(28953,16),
    to_signed(11272,16),
    to_signed(19005,16),
    to_signed(26708,16),
    to_signed(8934,16),
    to_signed(29220,16),
    to_signed(17893,16),
    to_signed(15717,16),
    to_signed(31339,16),
    to_signed(11048,16),
    to_signed(26601,16),
    to_signed(24287,16),
    to_signed(12755,16),
    to_signed(32767,16),
    to_signed(14651,16),
    to_signed(21945,16),
    to_signed(29204,16),
    to_signed(10982,16),
    to_signed(30816,16),
    to_signed(19035,16),
    to_signed(16403,16),
    to_signed(31567,16),
    to_signed(10819,16),
    to_signed(25915,16),
    to_signed(23145,16),
    to_signed(11159,16),
    to_signed(30719,16),
    to_signed(12155,16),
    to_signed(19005,16),
    to_signed(25824,16),
    to_signed(7168,16),
    to_signed(26574,16),
    to_signed(14373,16),
    to_signed(11327,16),
    to_signed(26087,16),
    to_signed(4942,16),
    to_signed(19652,16),
    to_signed(16505,16),
    to_signed(4153,16),
    to_signed(23359,16),
    to_signed(4453,16),
    to_signed(10973,16),
    to_signed(17475,16),
    to_signed(-1485,16),
    to_signed(17632,16),
    to_signed(5156,16),
    to_signed(1850,16),
    to_signed(16365,16),
    to_signed(-5008,16),
    to_signed(9489,16),
    to_signed(6146,16),
    to_signed(-6385,16),
    to_signed(12659,16),
    to_signed(-6393,16),
    to_signed(0,16),
    to_signed(6393,16),
    to_signed(-12659,16),
    to_signed(6385,16),
    to_signed(-6146,16),
    to_signed(-9489,16),
    to_signed(5008,16),
    to_signed(-16365,16),
    to_signed(-1850,16),
    to_signed(-5156,16),
    to_signed(-17632,16),
    to_signed(1485,16),
    to_signed(-17475,16),
    to_signed(-10973,16),
    to_signed(-4453,16),
    to_signed(-23359,16),
    to_signed(-4153,16),
    to_signed(-16505,16),
    to_signed(-19652,16),
    to_signed(-4942,16),
    to_signed(-26087,16),
    to_signed(-11327,16),
    to_signed(-14373,16),
    to_signed(-26574,16),
    to_signed(-7168,16),
    to_signed(-25824,16),
    to_signed(-19005,16),
    to_signed(-12155,16),
    to_signed(-30719,16),
    to_signed(-11159,16),
    to_signed(-23145,16),
    to_signed(-25915,16),
    to_signed(-10819,16),
    to_signed(-31567,16),
    to_signed(-16403,16),
    to_signed(-19035,16),
    to_signed(-30816,16),
    to_signed(-10982,16),
    to_signed(-29204,16),
    to_signed(-21945,16),
    to_signed(-14651,16),
    to_signed(-32767,16),
    to_signed(-12755,16),
    to_signed(-24287,16),
    to_signed(-26601,16),
    to_signed(-11048,16),
    to_signed(-31339,16),
    to_signed(-15717,16),
    to_signed(-17893,16),
    to_signed(-29220,16),
    to_signed(-8934,16),
    to_signed(-26708,16),
    to_signed(-19005,16),
    to_signed(-11272,16),
    to_signed(-28953,16),
    to_signed(-8514,16),
    to_signed(-19625,16),
    to_signed(-21526,16),
    to_signed(-5567,16),
    to_signed(-25462,16),
    to_signed(-9453,16),
    to_signed(-11253,16),
    to_signed(-22214,16),
    to_signed(-1574,16),
    to_signed(-19005,16),
    to_signed(-10973,16),
    to_signed(-2922,16),
    to_signed(-20301,16),
    to_signed(428,16),
    to_signed(-10408,16),
    to_signed(-12049,16),
    to_signed(4154,16),
    to_signed(-15512,16),
    to_signed(710,16),
    to_signed(-894,16),
    to_signed(-11676,16),
    to_signed(9127,16),
    to_signed(-8160,16),
    to_signed(0,16),
    to_signed(8160,16),
    to_signed(-9127,16),
    to_signed(11676,16),
    to_signed(894,16),
    to_signed(-710,16),
    to_signed(15512,16),
    to_signed(-4154,16),
    to_signed(12049,16),
    to_signed(10408,16),
    to_signed(-428,16),
    to_signed(20301,16),
    to_signed(2922,16),
    to_signed(10973,16),
    to_signed(19005,16),
    to_signed(1574,16),
    to_signed(22214,16),
    to_signed(11253,16),
    to_signed(9453,16),
    to_signed(25462,16),
    to_signed(5567,16),
    to_signed(21526,16),
    to_signed(19625,16),
    to_signed(8514,16),
    to_signed(28953,16),
    to_signed(11272,16),
    to_signed(19005,16),
    to_signed(26708,16),
    to_signed(8934,16),
    to_signed(29220,16),
    to_signed(17893,16),
    to_signed(15717,16),
    to_signed(31339,16),
    to_signed(11048,16),
    to_signed(26601,16),
    to_signed(24287,16),
    to_signed(12755,16),
    to_signed(32767,16),
    to_signed(14651,16),
    to_signed(21945,16),
    to_signed(29204,16),
    to_signed(10982,16),
    to_signed(30816,16),
    to_signed(19035,16),
    to_signed(16403,16),
    to_signed(31567,16),
    to_signed(10819,16),
    to_signed(25915,16),
    to_signed(23145,16),
    to_signed(11159,16),
    to_signed(30719,16),
    to_signed(12155,16),
    to_signed(19005,16),
    to_signed(25824,16),
    to_signed(7168,16),
    to_signed(26574,16),
    to_signed(14373,16),
    to_signed(11327,16),
    to_signed(26087,16),
    to_signed(4942,16),
    to_signed(19652,16),
    to_signed(16505,16),
    to_signed(4153,16),
    to_signed(23359,16),
    to_signed(4453,16),
    to_signed(10973,16),
    to_signed(17475,16),
    to_signed(-1485,16),
    to_signed(17632,16),
    to_signed(5156,16),
    to_signed(1850,16),
    to_signed(16365,16),
    to_signed(-5008,16),
    to_signed(9489,16),
    to_signed(6146,16),
    to_signed(-6385,16),
    to_signed(12659,16),
    to_signed(-6393,16),
    to_signed(0,16),
    to_signed(6393,16),
    to_signed(-12659,16),
    to_signed(6385,16),
    to_signed(-6146,16),
    to_signed(-9489,16),
    to_signed(5008,16),
    to_signed(-16365,16),
    to_signed(-1850,16),
    to_signed(-5156,16),
    to_signed(-17632,16),
    to_signed(1485,16),
    to_signed(-17475,16),
    to_signed(-10973,16),
    to_signed(-4453,16),
    to_signed(-23359,16),
    to_signed(-4153,16),
    to_signed(-16505,16),
    to_signed(-19652,16),
    to_signed(-4942,16),
    to_signed(-26087,16),
    to_signed(-11327,16),
    to_signed(-14373,16),
    to_signed(-26574,16),
    to_signed(-7168,16),
    to_signed(-25824,16),
    to_signed(-19005,16),
    to_signed(-12155,16),
    to_signed(-30719,16),
    to_signed(-11159,16),
    to_signed(-23145,16),
    to_signed(-25915,16),
    to_signed(-10819,16),
    to_signed(-31567,16),
    to_signed(-16403,16),
    to_signed(-19035,16),
    to_signed(-30816,16),
    to_signed(-10982,16),
    to_signed(-29204,16),
    to_signed(-21945,16),
    to_signed(-14651,16),
    to_signed(-32767,16),
    to_signed(-12755,16),
    to_signed(-24287,16),
    to_signed(-26601,16),
    to_signed(-11048,16),
    to_signed(-31339,16),
    to_signed(-15717,16),
    to_signed(-17893,16),
    to_signed(-29220,16),
    to_signed(-8934,16),
    to_signed(-26708,16),
    to_signed(-19005,16),
    to_signed(-11272,16),
    to_signed(-28953,16),
    to_signed(-8514,16),
    to_signed(-19625,16),
    to_signed(-21526,16),
    to_signed(-5567,16),
    to_signed(-25462,16),
    to_signed(-9453,16),
    to_signed(-11253,16),
    to_signed(-22214,16),
    to_signed(-1574,16),
    to_signed(-19005,16),
    to_signed(-10973,16),
    to_signed(-2922,16),
    to_signed(-20301,16),
    to_signed(428,16),
    to_signed(-10408,16),
    to_signed(-12049,16),
    to_signed(4154,16),
    to_signed(-15512,16),
    to_signed(710,16),
    to_signed(-894,16),
    to_signed(-11676,16),
    to_signed(9127,16),
    to_signed(-8160,16),
    to_signed(0,16),
    to_signed(8160,16),
    to_signed(-9127,16),
    to_signed(11676,16),
    to_signed(894,16),
    to_signed(-710,16),
    to_signed(15512,16),
    to_signed(-4154,16),
    to_signed(12049,16),
    to_signed(10408,16),
    to_signed(-428,16),
    to_signed(20301,16),
    to_signed(2922,16),
    to_signed(10973,16),
    to_signed(19005,16),
    to_signed(1574,16),
    to_signed(22214,16),
    to_signed(11253,16),
    to_signed(9453,16),
    to_signed(25462,16),
    to_signed(5567,16),
    to_signed(21526,16),
    to_signed(19625,16),
    to_signed(8514,16),
    to_signed(28953,16),
    to_signed(11272,16),
    to_signed(19005,16),
    to_signed(26708,16),
    to_signed(8934,16),
    to_signed(29220,16),
    to_signed(17893,16),
    to_signed(15717,16),
    to_signed(31339,16),
    to_signed(11048,16),
    to_signed(26601,16),
    to_signed(24287,16),
    to_signed(12755,16),
    to_signed(32767,16),
    to_signed(14651,16),
    to_signed(21945,16),
    to_signed(29204,16),
    to_signed(10982,16),
    to_signed(30816,16),
    to_signed(19035,16),
    to_signed(16403,16),
    to_signed(31567,16),
    to_signed(10819,16),
    to_signed(25915,16),
    to_signed(23145,16),
    to_signed(11159,16),
    to_signed(30719,16),
    to_signed(12155,16),
    to_signed(19005,16),
    to_signed(25824,16),
    to_signed(7168,16),
    to_signed(26574,16),
    to_signed(14373,16),
    to_signed(11327,16),
    to_signed(26087,16),
    to_signed(4942,16),
    to_signed(19652,16),
    to_signed(16505,16),
    to_signed(4153,16),
    to_signed(23359,16),
    to_signed(4453,16),
    to_signed(10973,16),
    to_signed(17475,16),
    to_signed(-1485,16),
    to_signed(17632,16),
    to_signed(5156,16),
    to_signed(1850,16),
    to_signed(16365,16),
    to_signed(-5008,16),
    to_signed(9489,16),
    to_signed(6146,16),
    to_signed(-6385,16),
    to_signed(12659,16),
    to_signed(-6393,16),
    to_signed(0,16),
    to_signed(6393,16),
    to_signed(-12659,16),
    to_signed(6385,16),
    to_signed(-6146,16),
    to_signed(-9489,16),
    to_signed(5008,16),
    to_signed(-16365,16),
    to_signed(-1850,16),
    to_signed(-5156,16),
    to_signed(-17632,16),
    to_signed(1485,16),
    to_signed(-17475,16),
    to_signed(-10973,16),
    to_signed(-4453,16),
    to_signed(-23359,16),
    to_signed(-4153,16),
    to_signed(-16505,16),
    to_signed(-19652,16),
    to_signed(-4942,16),
    to_signed(-26087,16),
    to_signed(-11327,16),
    to_signed(-14373,16),
    to_signed(-26574,16),
    to_signed(-7168,16),
    to_signed(-25824,16),
    to_signed(-19005,16),
    to_signed(-12155,16),
    to_signed(-30719,16),
    to_signed(-11159,16),
    to_signed(-23145,16),
    to_signed(-25915,16),
    to_signed(-10819,16),
    to_signed(-31567,16),
    to_signed(-16403,16),
    to_signed(-19035,16),
    to_signed(-30816,16),
    to_signed(-10982,16),
    to_signed(-29204,16),
    to_signed(-21945,16),
    to_signed(-14651,16),
    to_signed(-32767,16),
    to_signed(-12755,16),
    to_signed(-24287,16),
    to_signed(-26601,16),
    to_signed(-11048,16),
    to_signed(-31339,16),
    to_signed(-15717,16),
    to_signed(-17893,16),
    to_signed(-29220,16),
    to_signed(-8934,16),
    to_signed(-26708,16),
    to_signed(-19005,16),
    to_signed(-11272,16),
    to_signed(-28953,16),
    to_signed(-8514,16),
    to_signed(-19625,16),
    to_signed(-21526,16),
    to_signed(-5567,16),
    to_signed(-25462,16),
    to_signed(-9453,16),
    to_signed(-11253,16),
    to_signed(-22214,16),
    to_signed(-1574,16),
    to_signed(-19005,16),
    to_signed(-10973,16),
    to_signed(-2922,16),
    to_signed(-20301,16),
    to_signed(428,16),
    to_signed(-10408,16),
    to_signed(-12049,16),
    to_signed(4154,16),
    to_signed(-15512,16),
    to_signed(710,16),
    to_signed(-894,16),
    to_signed(-11676,16),
    to_signed(9127,16),
    to_signed(-8160,16),
    to_signed(0,16),
    to_signed(8160,16),
    to_signed(-9127,16),
    to_signed(11676,16),
    to_signed(894,16),
    to_signed(-710,16),
    to_signed(15512,16),
    to_signed(-4154,16),
    to_signed(12049,16),
    to_signed(10408,16),
    to_signed(-428,16),
    to_signed(20301,16),
    to_signed(2922,16),
    to_signed(10973,16),
    to_signed(19005,16),
    to_signed(1574,16),
    to_signed(22214,16),
    to_signed(11253,16),
    to_signed(9453,16),
    to_signed(25462,16),
    to_signed(5567,16),
    to_signed(21526,16),
    to_signed(19625,16),
    to_signed(8514,16),
    to_signed(28953,16),
    to_signed(11272,16),
    to_signed(19005,16),
    to_signed(26708,16),
    to_signed(8934,16),
    to_signed(29220,16),
    to_signed(17893,16),
    to_signed(15717,16),
    to_signed(31339,16),
    to_signed(11048,16),
    to_signed(26601,16),
    to_signed(24287,16),
    to_signed(12755,16),
    to_signed(32767,16),
    to_signed(14651,16),
    to_signed(21945,16),
    to_signed(29204,16),
    to_signed(10982,16),
    to_signed(30816,16),
    to_signed(19035,16),
    to_signed(16403,16),
    to_signed(31567,16),
    to_signed(10819,16),
    to_signed(25915,16),
    to_signed(23145,16),
    to_signed(11159,16),
    to_signed(30719,16),
    to_signed(12155,16),
    to_signed(19005,16),
    to_signed(25824,16),
    to_signed(7168,16),
    to_signed(26574,16),
    to_signed(14373,16),
    to_signed(11327,16),
    to_signed(26087,16),
    to_signed(4942,16),
    to_signed(19652,16),
    to_signed(16505,16),
    to_signed(4153,16),
    to_signed(23359,16),
    to_signed(4453,16),
    to_signed(10973,16),
    to_signed(17475,16),
    to_signed(-1485,16),
    to_signed(17632,16),
    to_signed(5156,16),
    to_signed(1850,16),
    to_signed(16365,16),
    to_signed(-5008,16),
    to_signed(9489,16),
    to_signed(6146,16),
    to_signed(-6385,16),
    to_signed(12659,16),
    to_signed(-6393,16),
    to_signed(0,16),
    to_signed(6393,16),
    to_signed(-12659,16),
    to_signed(6385,16),
    to_signed(-6146,16),
    to_signed(-9489,16),
    to_signed(5008,16),
    to_signed(-16365,16),
    to_signed(-1850,16),
    to_signed(-5156,16),
    to_signed(-17632,16),
    to_signed(1485,16),
    to_signed(-17475,16),
    to_signed(-10973,16),
    to_signed(-4453,16),
    to_signed(-23359,16),
    to_signed(-4153,16),
    to_signed(-16505,16),
    to_signed(-19652,16),
    to_signed(-4942,16),
    to_signed(-26087,16),
    to_signed(-11327,16),
    to_signed(-14373,16),
    to_signed(-26574,16),
    to_signed(-7168,16),
    to_signed(-25824,16),
    to_signed(-19005,16),
    to_signed(-12155,16),
    to_signed(-30719,16),
    to_signed(-11159,16),
    to_signed(-23145,16),
    to_signed(-25915,16),
    to_signed(-10819,16),
    to_signed(-31567,16),
    to_signed(-16403,16),
    to_signed(-19035,16),
    to_signed(-30816,16),
    to_signed(-10982,16),
    to_signed(-29204,16),
    to_signed(-21945,16),
    to_signed(-14651,16),
    to_signed(-32767,16),
    to_signed(-12755,16),
    to_signed(-24287,16),
    to_signed(-26601,16),
    to_signed(-11048,16),
    to_signed(-31339,16),
    to_signed(-15717,16),
    to_signed(-17893,16),
    to_signed(-29220,16),
    to_signed(-8934,16),
    to_signed(-26708,16),
    to_signed(-19005,16),
    to_signed(-11272,16),
    to_signed(-28953,16),
    to_signed(-8514,16),
    to_signed(-19625,16),
    to_signed(-21526,16),
    to_signed(-5567,16),
    to_signed(-25462,16),
    to_signed(-9453,16),
    to_signed(-11253,16),
    to_signed(-22214,16),
    to_signed(-1574,16),
    to_signed(-19005,16),
    to_signed(-10973,16),
    to_signed(-2922,16),
    to_signed(-20301,16),
    to_signed(428,16),
    to_signed(-10408,16),
    to_signed(-12049,16),
    to_signed(4154,16),
    to_signed(-15512,16),
    to_signed(710,16),
    to_signed(-894,16),
    to_signed(-11676,16),
    to_signed(9127,16),
    to_signed(-8160,16)
); 


begin

    -- Process for updating the filter with pipelined calculations
    process(clk, reset)
    variable index: integer:= 0; 
    begin
        if reset = '1' then
            -- Reset input and output registers to 0
            x_reg <= (others => (others => '0'));
            y_reg <= (others => (others => '0'));
            
            mul_x <= (others => (others => '0'));
            mul_y <= (others => (others => '0'));
            
            Sum_x <= (others => (others => '0'));
            Sum_y <= (others => (others => '0'));
            
            sample_valid_out <= '0';
            busy <= '0';
            state <= 0;
            index:=0; 
            
            --for debugging only
--            Flag <='1'; 
--            x_reg(0) <= to_signed(32767, 32); --signed(x_in);
        
        elsif rising_edge(clk) then
            case state is

                -- Initial stage: Load the input values and shift registers
                when 0 =>
                    if sample_validin_Sig = '1'  then
                       -- Shift input and output registers
                       x_in_Sig <= InputData(index);
                       x_reg(0) <= resize(signed(InputData(index)),32); --resize(signed(x_in),32); -- to_signed(32767, 16); --signed(x_in);
                       
                       index:= index+1; 
                       if(index = 1560) then 
                         index :=0; 
                       end if; 
                       
                       state <= 1;
                       busy <= '1';
                    end if;

                -- Stage 1: Multiply input values by coefficients
                when 1 =>
                
                    --Flag <='0'; 
                   
                    
                    for i in 0 to 6 loop
                        mul_x(i) <= x_reg(i) * b(i);  --8 bits * 16 bits  ==> need 24 bits
                    end loop;

                    -- Multiply previous output by feedback coefficients
                    for i in 1 to 6 loop
                       mul_y(i) <= y_reg(i) * a(i);  --8 bits * 16 bits  ==> need 24 bits
                    end loop;

                    state <= 2;

                -- Stage 2: Sum the multiplications
                when 2 =>
                    Sum_x(0) <= resize(mul_x(0) + mul_x(1),64);  
                    Sum_x(1) <= resize(mul_x(2) + mul_x(3),64);  
                    Sum_x(2) <= resize(mul_x(4) + mul_x(5),64);
                                                                 
                         
                    Sum_y(0) <= resize(mul_y(1) + mul_y(2),64);   
                    Sum_y(1) <= resize(mul_y(3) + mul_y(4),64); 
                    Sum_y(2) <= resize(mul_y(5) + mul_y(6),64);   

                    state <= 3;
                    
                 when 3 =>
                    Sum_x(3) <= resize(Sum_x(0) + Sum_x(1),64);    
                    Sum_x(4) <= resize(Sum_x(2) + mul_x(6),64);        
                                                                    
                    Sum_y(3) <= resize(Sum_y(0) + Sum_y(1),64);
                    
                    state <= 4; 
                    
                when 4 =>
                
                    Sum_x(5) <= resize(Sum_x(3) + Sum_x(4),64);             
                                                                             
                    Sum_y(4) <= resize(Sum_y(3) + Sum_y(2),64);               
                                                                            
                    state <= 5;
                    
                -- Stage 4: Reset output and prepare for next sample
                when 5 =>
  
                  OutputX <= Sum_x(5)- Sum_y(4);
                   
                   
                state <= 6;
                    
                when 6 => 
                    
                   Output <= resize(shift_right(OutputX,24),32);   --scale down by 2^24
                   
                   state <= 7;
                    
                   when 7 =>   
                   
                   --y_reg(1)<=  resize(Output,64);
                   y_reg(1)<=  Output;
                   
                     for i in 1 to 6 loop
                            x_reg(i) <= x_reg(i-1);
                        end loop;
              
                        for i in 2 to 6 loop
                            y_reg(i) <= y_reg(i-1);
                        end loop;
                    
                    sample_valid_out <= '1';
                    
                    state <= 8;

                    when 8 => 
                    
                    --for debugging only
                   -- x_reg(0) <= to_signed(0, 32); --signed(x_in);
                     
                    sample_valid_out <= '0';
                    busy <= '0';
                    state <= 0;
                 
                when others =>
                    state <= 0;
            end case;
        end if;
    end process;


 --   Output <= OutputX - OutputY; 

    -- Assign the output signal y[n] (output in Q0.16 format)
    iir_out <= std_logic_vector(output(15 downto 0));


-----------testing process-----------
--generate sample_valid_in ---
--syetm clock is 399.36
process(clk,reset)

begin
  if(reset='1') then
    clockcounter<=0;
    sample_validin_Sig<='0';
  elsif(rising_edge(clk)) then
    clockcounter <=clockcounter+1;
      if (clockcounter=64) then
          sample_validin_Sig <='1'; 
          clockcounter<=0; 
          else
          sample_validin_Sig <='0'; 
      end if;
    end if; 
end process;


sample_valid_in <= sample_validin_Sig; 


end Behavioral;
